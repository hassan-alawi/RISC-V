localparam NUM_INSTRUCTIONS = 5;